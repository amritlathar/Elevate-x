module full_subtractor (
    input A, B, Bin,  // A - B - Bin
    output Diff, Bout
);
    wire A_xor_B;
    xor (A_xor_B, A, B);      // Difference = A ^ B
    xor (Diff, A_xor_B, Bin); // Diff = (A ^ B) ^ Bin
    wire A_nand_B;
    nand (A_nand_B, A, B);
    wire not_A_xor_B, not_Bin;
    not (not_A_xor_B, A_xor_B);
    not (not_Bin, Bin);
    wire borrow1, borrow2;
    and (borrow1, not_A_xor_B, Bin);  // Borrow generated by Bin
    and (borrow2, A_nand_B, not_Bin); // Borrow generated by A and B
    or (Bout, borrow1, borrow2);  // Combine borrows
endmodule

module subtractor_3bit (
    input [2:0] A, B,     // Inputs to be subtracted (A - B)
    output [2:0] Diff,    // Difference
    output Bout           // Borrow out
);
    wire b1, b2;          // Internal borrow signals

    // Three full subtractors for 3-bit subtraction
    full_subtractor fs0 (A[0], B[0], 1'b0, Diff[0], b1);
    full_subtractor fs1 (A[1], B[1], b1, Diff[1], b2);
    full_subtractor fs2 (A[2], B[2], b2, Diff[2], Bout);
endmodule

module comparator_3bit (
    input [2:0] A, B,
    output A_less_B, A_equal_B, A_greater_B
);
    wire [2:0] A_xor_B;
    wire A_eq_0, A_eq_1, A_eq_2;

    // XOR to find where A and B differ
    xor (A_xor_B[0], A[0], B[0]);
    xor (A_xor_B[1], A[1], B[1]);
    xor (A_xor_B[2], A[2], B[2]);

    // A == B logic
    nor (A_eq_0, A_xor_B[0], A_xor_B[1], A_xor_B[2]);
    assign A_equal_B = A_eq_0;

    // A < B logic
    wire a2_b2, a1_b1, a0_b0;
    and (a2_b2, ~A[2], B[2]);  // A2 < B2
    and (a1_b1, ~A[1], B[1], ~A_xor_B[2]); // A1 < B1 when A2 == B2
    and (a0_b0, ~A[0], B[0], ~A_xor_B[1], ~A_xor_B[2]); // A0 < B0 when A1 == B1

    or (A_less_B, a2_b2, a1_b1, a0_b0);

    // A > B logic (A greater than B)
    assign A_greater_B = ~A_less_B & ~A_equal_B;
endmodule



module priority_controller (
    input [2:0] curr_floor_L1, curr_floor_L2,   // Current floors of Lift 1 and Lift 2
    input [2:0] dest_floor_L1, dest_floor_L2,   // Destination floors of Lift 1 and Lift 2
    input [2:0] req_floor,                      // Requested floor
    input req_direction,                        // Requested direction (1 = up, 0 = down)
    output [1:0] selected_lift                  // 00 = none, 01 = Lift 1, 10 = Lift 2
);

    wire [2:0] dist_L1, dist_L2;
    wire L1_less_L2, L1_equal_L2, L1_greater_L2;
    wire L1_moving_up, L2_moving_up, L1_moving_down, L2_moving_down;
    wire L1_prioritize, L2_prioritize;

    // Subtract distances using subtractor logic
    subtractor_3bit sub_L1 (.A(curr_floor_L1), .B(req_floor), .Diff(dist_L1), .Bout());
    subtractor_3bit sub_L2 (.A(curr_floor_L2), .B(req_floor), .Diff(dist_L2), .Bout());

    // Compare distances using comparator logic
    comparator_3bit comp_dist (.A(dist_L1), .B(dist_L2), .A_less_B(L1_less_L2), .A_equal_B(L1_equal_L2), .A_greater_B(L1_greater_L2));

    // Lift direction detection (moving up or down)
    wire L1_dir, L2_dir;
    wire not_req_direction, not_L1_moving_up, not_L2_moving_up;

    xor (L1_moving_up, curr_floor_L1[2], dest_floor_L1[2]); // XOR to detect lift direction
    xor (L2_moving_up, curr_floor_L2[2], dest_floor_L2[2]);

    not (L1_moving_down, L1_moving_up);
    not (L2_moving_down, L2_moving_up);

    // Prioritizing based on direction and proximity
    wire mux_L1_selected, mux_L2_selected;
    wire L1_less_L2_with_dir, L1_greater_L2_with_dir;

    and (L1_less_L2_with_dir, L1_less_L2, L1_moving_up);  // Prioritize Lift 1 if it's closer and moving up
    and (L1_greater_L2_with_dir, L1_greater_L2, L2_moving_up);  // Prioritize Lift 2 if it's closer and moving up

    or (mux_L1_selected, L1_less_L2_with_dir, L1_moving_down);
    or (mux_L2_selected, L1_greater_L2_with_dir, L2_moving_down);

    // Final lift selection logic
    assign selected_lift = (mux_L1_selected) ? 2'b01 : (mux_L2_selected ? 2'b10 : 2'b00);
endmodule

